library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fsm is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end fsm;

architecture rtl of fsm is

begin

end architecture;