library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SMDB is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end SMDB;

architecture rtl of SMDB is

begin

end architecture;