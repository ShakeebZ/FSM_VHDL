library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ControlUnit is
    port (
        clkCU : in std_logic;
        rstCU : in std_logic;
        hard_rstCU : in std_logic;
        instCU : in std_logic_vector(6 DOWNTO 0);
        toSegCU : out std_logic_vector(39 DOWNTO 0)
    );
end ControlUnit;

architecture rtl of ControlUnit is

begin

--PROCESS(rising_edge(clk))
--begin
toSegCU <= "0000000000000000000000000000000000000000" when (hard_rstCU = '1' OR instCU = "0000000" 
        OR (rstCU = '1' AND instCU(6) /= '1' AND instCU(5) /= '1')) ELSE
         "0000000000000000000000000000000000001010" when instCU = "0000001" ELSE --Program 1 Start
         "0000000000000000000000000000000101010001" when instCU = "0000010" ELSE
         "0000000000000000000000000010101000101011" when instCU = "0000011" ELSE
         "0000000000000000000001010100010101100000" when instCU = "0000100" ELSE
         "0000000000000000101010001010110000010110" when instCU = "0000101" ELSE
         "0000000000010101000101011000001011001010" when instCU = "0000110" ELSE
         "0000001010100010101100000101100101001110" when instCU = "0000111" ELSE
         "0101010001010110000010110010100111000000" when instCU = "0001000" ELSE
         "1000101011000001011001010011100000010100" when instCU = "0001001" ELSE
         "0101100000101100101001110000001010010101" when instCU = "0001010" ELSE
         "0000010110010100111000000101001010100101" when instCU = "0001011" ELSE
         "1011001010011100000010100101010010101111" when instCU = "0001100" ELSE
         "0101001110000001010010101001010111101111" when instCU = "0001101" ELSE
         "0111000000101001010100101011110111100101" when instCU = "0001110" ELSE
         "0000010100101010010101111011110010101111" when instCU = "0001111" ELSE
         "1010010101001010111101111001010111101101" when instCU = "0010000" ELSE
         "1010100101011110111100101011110110100000" when instCU = "0010001" ELSE
         "0010101111011110010101111011010000010010" when instCU = "0010010" ELSE
         "0111101111001010111101101000001001010000" when instCU = "0010011" ELSE
         "0111100101011110110100000100101000001111" when instCU = "0010100" ELSE
         "0010101111011010000010010100000111100000" when instCU = "0010101" ELSE
         "0111101101000001001010000011110000000000" when instCU = "0010110" ELSE
         "0110100000100101000001111000000000001111" when instCU = "0010111" ELSE
         "0000010010100000111100000000000111110000" when instCU = "0011000" ELSE
         "1001010000011110000000000011111000000000" when instCU = "0011001" ELSE
         "1000001111000000000001111100000000000000" when instCU = "0011010" ELSE
         "0111100000000000111110000000000000000000" when instCU = "0011011" ELSE
         "0000000000011111000000000000000000000000" when instCU = "0011100" ELSE
         "0000001111100000000000000000000000000000" when instCU = "0011101" ELSE
         "0111110000000000000000000000000000000000" when instCU = "0011110" ELSE
         "1000000000000000000000000000000000000000" when instCU = "0011111" ELSE -- Program 1 End
         "0000000000000000000000000000000000000111" when instCU = "0100000" ELSE -- Program 2 Start
         "0000000000000000000000000000000011101001" when instCU = "0100001" ELSE
         "0000000000000000000000111010010100111000" when instCU = "0100010" ELSE
         "0000000000000000011101001010011100011000" when instCU = "0100011" ELSE
         "0000000000001110100101001110001100000000" when instCU = "0100100" ELSE
         "0000000111010010100111000110000000000000" when instCU = "0100101" ELSE
         "0011101001010011100011000000000000000000" when instCU = "0100110" ELSE
         "0100101001110001100000000000000000000000" when instCU = "0100111" ELSE
         "0100111000110000000000000000000000000000" when instCU = "0101000" ELSE
         "1100011000000000000000000000000000000000" when instCU = "0101001" ELSE
         "1100000000000000000000000000000000000000" when instCU = "0101010" ELSE -- Program 2 End
         "0100000000000000000000000000000000000000" when instCU = "0101011" ELSE -- Program 3 Start
         "0100101000000000000000000000000000000000" when instCU = "0101100" ELSE
         "0100101001010000000000000000000000000000" when instCU = "0101101" ELSE
         "1010101001010010100000000000000000000000" when instCU = "0101110" ELSE
         "0000010101010010100101000000000000000000" when instCU = "0101111" ELSE
         "0000000000101010100101001010000000000000" when instCU = "0110000" ELSE
         "0000000000000001010101001010010100000000" when instCU = "0110001" ELSE
         "0000000000000000000010101010010100101000" when instCU = "0110010" ELSE
         "0000000000000000000000000101010100101001" when instCU = "0110011" ELSE
         "0000000000000000000000000000001010101001" when instCU = "0110100" ELSE
         "0000000000000000000000000000000000010101" when instCU = "0110101" ELSE -- Program 3 End
         "0000000000000000000000000000000000000001" when instCU = "1100000" ELSE -- Program 4 Start
         "0000000000000000000000000000000000000100" when instCU = "1100001" ELSE
         "0000000000000000000000000000000000000010" when instCU = "1100010" ELSE
         "0000000000000000000000000000000000000110" when instCU = "1100011" ELSE
         "0000000000000000000000000000000000000110" when instCU = "1100100" ELSE
         "0000000000000000000000000000000000000011" when instCU = "1100101" ELSE
         "0000000000000000000000000000000000010111" when instCU = "1100110" ELSE
         "0000000000000000000000000000000000000101" when instCU = "1100111" ELSE
         "0000000000000000000000000000000000000110" when instCU = "1101000" ELSE
         "0000000000000000000000000000000000100000" when instCU = "1101001" ELSE
         "0000000000000000000000000000000010000000" when instCU = "1101010" ELSE
         "0000000000000000000000000000000001000000" when instCU = "1101011" ELSE
         "0000000000000000000000000000000011000000" when instCU = "1101100" ELSE 
         "0000000000000000000000000000000000000110" when instCU = "1101101" ELSE
         "0000000000000000000000000000000001100000" when instCU = "1101110" ELSE
         "0000000000000000000000000000001011100000" when instCU = "1101111" ELSE
         "0000000000000000000000000000000010100000" when instCU = "1110000" ELSE
         "0000000000000000000000000000000000000110" when instCU = "1110001" ELSE -- Program 4 End
         "0000000000011000101000101110000000000000" when instCU = "1110010" ELSE -- Error Message
         "0000000000000000000000000000000000000000";


--END PROCESS;

end architecture;