library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ToneGenerator is
    port (
        clkTG : in std_logic;
        instTG : in std_logic_vector(6 DOWNTO 0);
        AUD_ADCDAT
    );
end ToneGenerator;

architecture rtl of ToneGenerator is

begin

end architecture;